module some_module (
    input wire a,
    input wire b,
    output wire z
);

assign z = a && b;

endmodule
